<?xml version="1.0" encoding="UTF-8"?>
<svg xmlns="http://www.w3.org/2000/svg" version="1.1" width="100" height="100" viewBox="0 0 100 100"><rect x="0" y="0" width="100" height="100" fill="#ffffff"/><g transform="scale(4.762)"><g transform="translate(0,0)"><path fill-rule="evenodd" d="M9 0L9 1L8 1L8 3L9 3L9 4L8 4L8 8L6 8L6 9L4 9L4 8L3 8L3 9L2 9L2 8L0 8L0 9L1 9L1 10L0 10L0 13L1 13L1 12L2 12L2 13L5 13L5 12L6 12L6 13L8 13L8 15L10 15L10 16L11 16L11 18L9 18L9 17L8 17L8 18L9 18L9 19L8 19L8 21L13 21L13 20L16 20L16 21L17 21L17 20L18 20L18 19L19 19L19 18L20 18L20 19L21 19L21 15L20 15L20 14L21 14L21 13L20 13L20 12L21 12L21 9L20 9L20 8L18 8L18 9L17 9L17 8L14 8L14 10L12 10L12 11L11 11L11 12L12 12L12 13L11 13L11 14L12 14L12 13L13 13L13 12L12 12L12 11L14 11L14 10L16 10L16 9L17 9L17 10L18 10L18 11L19 11L19 13L18 13L18 15L17 15L17 14L16 14L16 16L17 16L17 17L16 17L16 19L13 19L13 18L12 18L12 16L14 16L14 17L15 17L15 16L14 16L14 14L13 14L13 15L10 15L10 13L9 13L9 12L10 12L10 10L11 10L11 8L13 8L13 4L12 4L12 3L13 3L13 2L12 2L12 1L13 1L13 0L11 0L11 2L12 2L12 3L11 3L11 4L12 4L12 5L11 5L11 6L10 6L10 7L9 7L9 4L10 4L10 0ZM11 6L11 7L12 7L12 6ZM8 8L8 9L9 9L9 10L7 10L7 9L6 9L6 10L5 10L5 11L6 11L6 12L7 12L7 11L9 11L9 10L10 10L10 9L9 9L9 8ZM3 9L3 10L4 10L4 9ZM18 9L18 10L19 10L19 11L20 11L20 9ZM1 10L1 11L2 11L2 12L3 12L3 11L2 11L2 10ZM6 10L6 11L7 11L7 10ZM15 11L15 12L14 12L14 13L17 13L17 12L16 12L16 11ZM19 13L19 14L20 14L20 13ZM18 15L18 17L17 17L17 18L19 18L19 17L20 17L20 15ZM11 18L11 19L9 19L9 20L13 20L13 19L12 19L12 18ZM16 19L16 20L17 20L17 19ZM19 20L19 21L20 21L20 20ZM0 0L0 7L7 7L7 0ZM1 1L1 6L6 6L6 1ZM2 2L2 5L5 5L5 2ZM14 0L14 7L21 7L21 0ZM15 1L15 6L20 6L20 1ZM16 2L16 5L19 5L19 2ZM0 14L0 21L7 21L7 14ZM1 15L1 20L6 20L6 15ZM2 16L2 19L5 19L5 16Z" fill="#000000"/></g></g></svg>
